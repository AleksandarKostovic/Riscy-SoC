`ifdefine OPCODES
`define OPCODES

`define INSTR_LUI     64'b???????_?????_?????_???_?????_0110111 /* LUI */
`define INSTR_AUIPC   64'b???????_?????_?????_???_?????_0010111 /* AUIPC */
`define INSTR_JAL     64'b???????_?????_?????_???_?????_1101111 /* JAL */
`define INSTR_JALR    64'b???????_?????_?????_000_?????_1100111 /* JALR */
`define INSTR_BEQ     64'b???????_?????_?????_000_?????_1100011 /* BRANCH */
`define INSTR_BNE     64'b???????_?????_?????_001_?????_1100011
`define INSTR_BLT     64'b???????_?????_?????_100_?????_1100011
`define INSTR_BGE     64'b???????_?????_?????_101_?????_1100011
`define INSTR_BLTU    64'b???????_?????_?????_110_?????_1100011
`define INSTR_BGEU    64'b???????_?????_?????_111_?????_1100011
`define INSTR_LB      64'b???????_?????_?????_000_?????_0000011 /* LOAD */
`define INSTR_LH      64'b???????_?????_?????_001_?????_0000011
`define INSTR_LW      64'b???????_?????_?????_010_?????_0000011
`define INSTR_LBU     64'b???????_?????_?????_100_?????_0000011
`define INSTR_LHU     64'b???????_?????_?????_101_?????_0000011
`define INSTR_SB      64'b???????_?????_?????_000_?????_0100011 /* STORE */
`define INSTR_SH      64'b???????_?????_?????_001_?????_0100011
`define INSTR_SW      64'b???????_?????_?????_010_?????_0100011
`define INSTR_ADDI    64'b???????_?????_?????_000_?????_0010011 /* OP-IMM */
`define INSTR_SLTI    64'b???????_?????_?????_010_?????_0010011
`define INSTR_SLTIU   64'b???????_?????_?????_011_?????_0010011
`define INSTR_XORI    64'b???????_?????_?????_100_?????_0010011
`define INSTR_ORI     64'b???????_?????_?????_110_?????_0010011
`define INSTR_ANDI    64'b???????_?????_?????_111_?????_0010011
`define INSTR_SLLI    64'b0000000_?????_?????_001_?????_0010011
`define INSTR_SRLI    64'b0000000_?????_?????_101_?????_0010011
`define INSTR_SRAI    64'b0100000_?????_?????_101_?????_0010011
`define INSTR_ADD     64'b0000000_?????_?????_000_?????_0110011 /* OP */
`define INSTR_SUB     64'b0100000_?????_?????_000_?????_0110011
`define INSTR_SLL     64'b0000000_?????_?????_001_?????_0110011
`define INSTR_SLT     64'b0000000_?????_?????_010_?????_0110011
`define INSTR_SLTU    64'b0000000_?????_?????_011_?????_0110011
`define INSTR_XOR     64'b0000000_?????_?????_100_?????_0110011
`define INSTR_SRL     64'b0000000_?????_?????_101_?????_0110011
`define INSTR_SRA     64'b0100000_?????_?????_101_?????_0110011
`define INSTR_OR      64'b0000000_?????_?????_110_?????_0110011
`define INSTR_AND     64'b0000000_?????_?????_111_?????_0110011
`define INSTR_FENCE   64'b???????_?????_?????_000_?????_0001111 /* MISC-MEM */
`define INSTR_FENCE_I 64'b???????_?????_?????_001_?????_0001111
`define INSTR_ECALL   64'b0000000_00000_00000_000_00000_1110011 /* SYSTEM */
`define INSTR_EBREAK  64'b0000000_00001_00000_000_00000_1110011
`define INSTR_MRET    64'b0011000_00010_00000_000_00000_1110011
`define INSTR_WFI     64'b0001000_00101_00000_000_00000_1110011
`define INSTR_CSRRW   64'b???????_?????_?????_001_?????_1110011
`define INSTR_CSRRS   64'b???????_?????_?????_010_?????_1110011
`define INSTR_CSRRC   64'b???????_?????_?????_011_?????_1110011
`define INSTR_CSRRWI  64'b???????_?????_?????_101_?????_1110011
`define INSTR_CSRRSI  64'b???????_?????_?????_110_?????_1110011
`define INSTR_CSRRCI  64'b???????_?????_?????_111_?????_1110011

`define INSTR_NOP     64'bxxxxxxx_xxxxx_00000_xxx_00000_0010011

`define OPCODE_JAL    7'b1101111
`define OPCODE_BRANCH 7'b1100011

`endif
