`define beg
`define bne
`define blt
`define bge
`define bltu
`define bgeu
`define jalr
`define jal
`define lui
`define auipc
`define addi
`define slli
`define slti 
`define sltiu 
`define xori 
`define srli
`define srai
`define ori
`define andi
`define add 
`define sub
`define sll
`define slt
`define sltu 
`define xor
`define srl 
`define sra 
`define or
`define and
`define addiw
`define slliw
`define srliw 
`define sraiw
`define addw
`define subw
`define sllw 
`define srlw
`define sraw
`define lb 
`define lh
`define lw
`define ld
`define lbu
`define lhu
`define lwu
`define sb
`define sh
`define sw
`define sd
`define fence
`define fence.i
`define mul
`define mulh
`define mulhsu
`define mulhu
`define div
`define divu
`define rem
`define remu 
`define mulw
`define divw
`define divuw
`define remw
`define remuw 
//to do:RVA and SYSTEM
