//ram
